library verilog;
use verilog.vl_types.all;
entity TestBench is
end TestBench;
